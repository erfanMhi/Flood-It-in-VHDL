----------------------------------------------------------------------------------
-- Moving Square Demonstration 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use ieee.numeric_std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

LIBRARY work;
use work.Graphic_Lab.all;
entity Board is
  port ( CLK_50MHz		: in std_logic;
			RESET				: in std_logic;
			ColorOut			: out std_logic_vector(11 downto 0); -- RED & GREEN & BLUE
			SQUAREWIDTH		: in std_logic_vector(7 downto 0);
			ScanlineX		: in std_logic_vector(10 downto 0);
			ScanlineY		: in std_logic_vector(10 downto 0)
  );
end Board;

architecture Behavioral of Board is
  
  shared variable ColorOutput: std_logic_vector(11 downto 0);
  
  signal column_width: std_logic_vector(9 downto 0) := "0000000001";
  signal row_width: std_logic_vector(9 downto 0) := "0000000001";
  
  signal food_size: std_logic_vector(10 downto 0) := "00000010110";
  signal food_inc: boolean:= false;
  
  signal SquareX: std_logic_vector(9 downto 0) := "0000001110";  
  signal SquareY: std_logic_vector(9 downto 0) := "0000010111";  
  signal SquareXMoveDir, SquareYMoveDir: std_logic := '0';
  --constant SquareWidth: std_logic_vector(4 downto 0) := "11001";
  constant SquareXmin: std_logic_vector(9 downto 0) := "0000000001";
  signal SquareXmax: std_logic_vector(9 downto 0); -- := "1010000000"-SquareWidth;
  constant SquareYmin: std_logic_vector(9 downto 0) := "0000000001";
  signal SquareYmax: std_logic_vector(9 downto 0); -- := "0111100000"-SquareWidth;
  signal ColorSelect: std_logic_vector(2 downto 0) := "001";
  signal Prescaler: std_logic_vector(40 downto 0) := (others => '0');

begin

	PrescalerCounter: process(CLK_50Mhz, RESET)
	begin
		if RESET = '1' then
			Prescaler <= (others => '0');
			SquareX <= "0111000101";
			SquareY <= "0001100010";
			SquareXMoveDir <= '0';
			SquareYMoveDir <= '0';
			ColorSelect <= "001";
		elsif rising_edge(CLK_50Mhz) then
			Prescaler <= Prescaler + 1;	 
			if Prescaler = "0000000000000000000100000000000000000000" then  -- Activated every 0,002 sec (2 msec)
				Prescaler <= (others => '0');
				if food_size = "00000010110" then
					food_inc <= false;
				elsif food_size = "00000000001" then
					food_inc <= true;
				end if;
				if food_inc = true then
					food_size <= food_size +1;
				else
					food_size <= food_size -1;
				end if;
			end if;
		end if;
	end process PrescalerCounter;
	
	color_painter: process(ScanlineX, ScanlineY)
	begin
		if (ScanlineX < std_logic_vector(to_unsigned(213, 10))) and
		(ScanlineX > std_logic_vector(to_unsigned(0, 10))) and
		(ScanlineY > std_logic_vector(to_unsigned(50, 10))) and
		(ScanlineY < std_logic_vector(to_unsigned(60, 10))) then
			ColorOutput := "111111000000";
		else  
			ColorOutput := "111111111111";
		end if;
		
		-- left arrow
		Coloroutput := draw_line(std_logic_vector(to_unsigned(300, 11)), std_logic_vector(to_unsigned(455, 11)), std_logic_vector(to_unsigned(330, 11)), std_logic_vector(to_unsigned(455, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(300, 11)), std_logic_vector(to_unsigned(455, 11)), std_logic_vector(to_unsigned(310, 11)), std_logic_vector(to_unsigned(445, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(300, 11)), std_logic_vector(to_unsigned(455, 11)), std_logic_vector(to_unsigned(310, 11)), std_logic_vector(to_unsigned(465, 11)), ScanlineX, ScanlineY);
		
		-- up arrow
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(335, 11)), std_logic_vector(to_unsigned(440, 11)), std_logic_vector(to_unsigned(335, 11)), std_logic_vector(to_unsigned(470, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(335, 11)), std_logic_vector(to_unsigned(440, 11)), std_logic_vector(to_unsigned(345, 11)), std_logic_vector(to_unsigned(450, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(335, 11)), std_logic_vector(to_unsigned(440, 11)), std_logic_vector(to_unsigned(325, 11)), std_logic_vector(to_unsigned(450, 11)), ScanlineX, ScanlineY);
		
		-- down arrow
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(355, 11)), std_logic_vector(to_unsigned(460, 11)), std_logic_vector(to_unsigned(345, 11)), std_logic_vector(to_unsigned(470, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(335, 11)), std_logic_vector(to_unsigned(460, 11)), std_logic_vector(to_unsigned(345, 11)), std_logic_vector(to_unsigned(470, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(345, 11)), std_logic_vector(to_unsigned(440, 11)), std_logic_vector(to_unsigned(345, 11)), std_logic_vector(to_unsigned(470, 11)), ScanlineX, ScanlineY);
		
		-- right arrow
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(380, 11)), std_logic_vector(to_unsigned(455, 11)), std_logic_vector(to_unsigned(350, 11)), std_logic_vector(to_unsigned(455, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(380, 11)), std_logic_vector(to_unsigned(455, 11)), std_logic_vector(to_unsigned(370, 11)), std_logic_vector(to_unsigned(465, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(380, 11)), std_logic_vector(to_unsigned(455, 11)), std_logic_vector(to_unsigned(370, 11)), std_logic_vector(to_unsigned(445, 11)), ScanlineX, ScanlineY);
		
		-- rectangle
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(80, 11)), std_logic_vector(to_unsigned(50, 11)), std_logic_vector(to_unsigned(600, 11)), std_logic_vector(to_unsigned(50, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(80, 11)), std_logic_vector(to_unsigned(50, 11)), std_logic_vector(to_unsigned(80, 11)), std_logic_vector(to_unsigned(430, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(600, 11)), std_logic_vector(to_unsigned(430, 11)), std_logic_vector(to_unsigned(80, 11)), std_logic_vector(to_unsigned(430, 11)), ScanlineX, ScanlineY);
		Coloroutput := Coloroutput and draw_line(std_logic_vector(to_unsigned(600, 11)), std_logic_vector(to_unsigned(430, 11)), std_logic_vector(to_unsigned(600, 11)), std_logic_vector(to_unsigned(50, 11)), ScanlineX, ScanlineY);
	
		-- colored cells
		ColorOutput :=	Coloroutput and colorize_cell("00000101111", "00000100110", ScanlineX, ScanlineY);
		ColorOutput :=	Coloroutput and colorize_cell("00000101110", "00000100110", ScanlineX, ScanlineY);
		ColorOutput :=	Coloroutput and colorize_cell("00000101110", "00000100111", ScanlineX, ScanlineY);
		ColorOutput :=	Coloroutput and colorize_cell("00000101110", "00000101000", ScanlineX, ScanlineY);
		--ColorOutput :=	Coloroutput and colorize_cell("00000100110", "00000010110", ScanlineX, ScanlineY);
		ColorOutput :=	Coloroutput and draw_circle("00000100110", "00000010110", food_size, ScanlineX, ScanlineY);
	end process;
	ColorOut <= ColorOutput;
	
	SquareXmax <= "1010000000"-SquareWidth; -- (640 - SquareWidth)
	SquareYmax <= "0111100000"-SquareWidth;	-- (480 - SquareWidth)
	
end Behavioral;

